// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by osboxes on Thu 20 Feb 01:56:03 EST 2020
//
// cmd:    swerv -snapshot=pynqz2 -ret_stack_size=8 -iccm_enable=0 dccm_enable=0 -fpga_optimize = 1 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG CKLNQD12BWP35P140
`define PHYSICAL 1
